module and_2(out, in_1, in_2);

output out;
input in_1, in_2;
assign out = in_1 & in_2;

endmodule
