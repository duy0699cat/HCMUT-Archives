module invert 
(
 input in,
 output out
 );
 
 assign out = ~in;
 
 endmodule 